module fulladd (  input [3:0] a,
                  input [3:0] b,
                output [3:0] sum);

   assign {sum} = a + b;
endmodule
